library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- This package is designed to define some constant used in the project.
package header is
    constant MEM_BITS               : INTEGER := 16;                                -- number of bits per word
    constant ADDR_BITS              : INTEGER := 8;                                 -- number of bits per address in memory
    -- TODO: set ENTRIES to be equal to 2^32
    constant ENTRIES                : INTEGER := 2 ** ADDR_BITS;                    -- number of entries
    -- TODO: set PCDelta to be equal to 32/MEM_BITS
    constant PCDelta                : STD_LOGIC_VECTOR(31 downto 0) := x"00000002"; -- number of PC added in each cycle

    constant OP_RType               : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"0";
    constant OP_ADDI                : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"1";
--  constant OP_SUB                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"0";
    constant OP_SUBI                : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"2";
--  constant OP_AND                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"0";
    constant OP_ANDI                : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"3";
--  constant OP_OR                  : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"0";
--  constant OP_NOR                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"0";
    constant OP_ORI                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"4";
    constant OP_SHR                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"5";
    constant OP_SHL                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"6";
        
    constant OP_LW                  : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"7";
    constant OP_SW                  : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"8";
    constant OP_BLT                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"9";
    constant OP_BEQ                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"A";
    constant OP_BNE                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"B";
    constant OP_JMP                 : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"C";

    constant OP_HAL                 : STD_LOGIC_VECTOR(5 downto 0) := "11" & x"F";
            
    constant FUNC_ADD               : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"1";
    constant FUNC_SUB               : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"3";
    constant FUNC_AND               : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"5";
    constant FUNC_OR                : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"7";
    constant FUNC_NOR               : STD_LOGIC_VECTOR(5 downto 0) := "00" & x"9";
            
    constant ALU_ADD                : STD_LOGIC_VECTOR(3 downto 0) := x"0";
    constant ALU_SUB                : STD_LOGIC_VECTOR(3 downto 0) := x"1";
    constant ALU_AND                : STD_LOGIC_VECTOR(3 downto 0) := x"2";
    constant ALU_OR                 : STD_LOGIC_VECTOR(3 downto 0) := x"3";
    constant ALU_NOR                : STD_LOGIC_VECTOR(3 downto 0) := x"4";
    constant ALU_SHR                : STD_LOGIC_VECTOR(3 downto 0) := x"5";
    -- constant ALU_SHL             : STD_LOGIC_VECTOR(3 downto 0) := x"6";
    constant ALU_BLT                : STD_LOGIC_VECTOR(3 downto 0) := x"7";
    constant ALU_BEQ                : STD_LOGIC_VECTOR(3 downto 0) := x"8";
    constant ALU_BNE                : STD_LOGIC_VECTOR(3 downto 0) := x"9";
    constant ALU_XOR                : STD_LOGIC_VECTOR(3 downto 0) := x"a";
    constant ALU_NDEF               : STD_LOGIC_VECTOR(3 downto 0) := x"f";

    type mem is array (0 to ENTRIES - 1) of STD_LOGIC_VECTOR(MEM_BITS - 1 downto 0);
    -- RC5 encryption
    constant instr_enc : mem := (
        -- initialize part
        -- R0 stores zero
        -- initialize R0 to be 0
        "0000000000000000","0000000000000011",          -- SUB R0, R0, R0
        -- R1 stores the input A
        "0001110000000001","0000000000110100",          -- LW R1 52(R0)
        -- R2 stores the input B
        "0001110000000010","0000000000110110",          -- LW R2 54(R0)
        -- R3 stores i
        -- initialize R3 to be 0
        "0000000001100011","0001100000000011",          -- SUB R3, R3, R3
        -- R6 stores S[0]
        "0001110000000110","0000000000000000",          -- LW R6, 0(R0)
        -- R7 stores S[1]
        "0001110000000111","0000000000000010",          -- LW R7, 2(R0)
        -- R8 stores intermediate A
        -- A = A + S[0]
        "0000000000100110","0100000000000001",          -- ADD R8, R1, R6
        -- R9 stores intermediate B
        -- B = B + S[1]
        "0000000001000111","0100100000000001",          -- ADD R9, R2, R7
        -- R10 stores 12
        "0000010000001010","0000000000001100",          -- ADDI R10, R0, 12
        
        -- encryption loop begin
        -- R3 = R3 + 1
        "0000010001100011","0000000000000001",          -- ADDI R3, R3, 1
        -- R4 stores 2*i
        "0000000001100011","0010000000000001",          -- ADD R4, R3, R3
        -- R5 stores 2*i+1
        "0000010010000101","0000000000000001",          -- ADDI R5, R4, 1
        -- R4 and R5 multiplied by 2 because 16-bit addressable
        "0000000010000100","0010000000000001",          -- ADD R4, R4, R4
        "0000000010100101","0010100000000001",          -- ADD R5, R5, R5
        -- R6 stores S[2*i]
        "0001110010000110","0000000000000000",          -- LW R6, 0(R4)
        -- R7 stores S[2*i+1]
        "0001110010100111","0000000000000000",          -- LW R7, 0(R5)

        -- A = A xor B
        -- R11 stores A nor B
        "0000000100001001","0101100000001001",          -- NOR R11, R8, R9
        -- R12 stores A and B
        "0000000100001001","0110000000000101",          -- AND R12, R8, R9
        -- A = A xor B = (A nor B) nor (A and B) 
        "0000000101101100","0100000000001001",          -- NOR R8, R11, R12

        -- A = A <<< B
        -- initialize R11 with A
        "0000010100001011","0000000000000000",          -- ADDI R11, R8, 0
        -- R13 stores B[4:0] - 32
        "0000110100101101","0000000000011111",          -- ANDI R13, R9, 31
        "0000100110101101","0000000000100000",          -- SUBI R13, R13, 32
        -- R11 loop begin
        "0010100110100000","0000000000000011",          -- BEQ R13, R0, 3
        -- R11 stores B[4:0] MSBs of A
        "0001010101101011","0000000000000001",          -- SHR R11, R11, 1
        -- R13 = R13 + 1
        "0000010110101101","0000000000000001",          -- ADDI R13, R13, 1
        -- R11 loop while R13 < 0
        "0010110110100000","1111111111111101",          -- BNE R13, R0, -3
        -- initialize R12 with A
        "0000010100001100","0000000000000000",          -- ADDI R12, R8, 0
        -- R13 stores B[4:0]
        "0000110100101101","0000000000011111",          -- ANDI R13, R9, 31
        -- R12 loop begin
        "0010100110100000","0000000000000011",          -- BEQ R13, R0, 3
        -- R12 stores A shifted by B[4:0] bits left
        "0000000110001100","0110000000000001",          -- ADD R12, R12, R12
        -- R13 = R13 - 1
        "0000100110101101","0000000000000001",          -- SUBI R13, R13, 1
        -- R12 loop while R13 > 0
        "0010110110100000","1111111111111101",          -- BNE R13, R0, -3
        -- A = R11 or R12
        "0000000101101100","0100000000000111",          -- OR R8, R11, R12

        -- A = A + S[2*i]
        "0000000100000110","0100000000000001",          -- ADD R8, R8, R6

        -- B = B xor A
        -- R11 stores B nor A
        "0000000100101000","0101100000001001",          -- NOR R11, R9, R8
        -- R12 stores B and A
        "0000000100101000","0110000000000101",          -- AND R12, R9, R8
        -- B = B xor A = (B nor A) nor (B and A) 
        "0000000101101100","0100100000001001",          -- NOR R9, R11, R12

        -- B = B <<< A
        -- initialize R11 with B
        "0000010100101011","0000000000000000",          -- ADDI R11, R9, 0
        -- R13 stores A[4:0] - 32
        "0000110100001101","0000000000011111",          -- ANDI R13, R8, 31
        "0000100110101101","0000000000100000",          -- SUBI R13, R13, 32
        -- R11 loop begin
        "0010100110100000","0000000000000011",          -- BEQ R13, R0, 3
        -- R11 stores A[4:0] MSBs of B
        "0001010101101011","0000000000000001",          -- SHR R11, R11, 1
        -- R13 = R13 + 1
        "0000010110101101","0000000000000001",          -- ADDI R13, R13, 1
        -- R11 loop while R13 < 0
        "0010110110100000","1111111111111101",          -- BNE R13, R0, -3
        -- initialize R12 with B
        "0000010100101100","0000000000000000",          -- ADDI R12, R9, 0
        -- R13 stores A[4:0]
        "0000110100001101","0000000000011111",          -- ANDI R13, R8, 31
        -- R12 loop begin
        "0010100110100000","0000000000000011",          -- BEQ R13, R0, 3
        -- R12 stores B shifted by A[4:0] bits left
        "0000000110001100","0110000000000001",          -- ADD R12, R12, R12
        -- R13 = R13 - 1
        "0000100110101101","0000000000000001",          -- SUBI R13, R13, 1
        -- R12 loop while R13 > 0
        "0010110110100000","1111111111111101",          -- BNE R13, R0, -3
        -- B = R11 or R12
        "0000000101101100","0100100000000111",          -- OR R9, R11, R12

        -- B = B + S[2*i+1]
        "0000000100100111","0100100000000001",          -- ADD R9, R9, R7
        
        -- encryption loop while i < 12
        "0010010001101010","1111111111010100",          -- BLT R3, R10, -44

        -- store encrypted A to Mem[56]
        "0010000000001000","0000000000111000",          -- SW R8, 56(R0)

        -- store encrypted B to Mem[58]
        "0010000000001001","0000000000111010",          -- SW R9, 58(R0)

        -- halt
        "1111110000000000","0000000000000000",          -- HAL
        others => x"0000"
    );

    -- RC5 deryption
    constant instr_dec : mem := (
        -- initialize part
        -- initialize R0 to 0
        "0000000000000000", "0000000000000011",         -- SUB R0, R0, R0
        -- R3 stores 13 
        "0000010000000011", "0000000000001101",         -- ADDI R3, R0, 13
        -- load A 
        "0001110000001000", "0000000000110100",         -- LW R8, 52(R0)
        -- load B 
        "0001110000001001", "0000000000110110",         -- LW R9, 54(R0)
        -- set R1 as 1 
        "0000010000000001", "0000000000000001",         -- ADDI R1, R0, 1
 
        -- decryption loop begins
        -- R3 = R3 -1 
        "0000100001100011", "0000000000000001",         -- SUBI R3, R3, 1
        -- R4 stores 2*i 
        "0000000001100011", "0010000000000001",         -- ADD R4, R3, R3
        -- R5 stores 2*i+1 
        "0000010010000101", "0000000000000001",         -- ADDI R5, R4, 1 
 
        -- R4 and R5 multiplied by 2 because 16-bit addressable
        "0000000010000100", "0010000000000001",         -- ADD R4, R4, R4
        "0000000010100101", "0010100000000001",         -- ADD R5, R5, R5
        -- R6 stores S[2*i] 
        "0001110010000110", "0000000000000000",         -- LW R6, 0(R4)
        -- R7 stores S[2*i+1]
        "0001110010100111", "0000000000000000",         -- LW R7, 0(R5)
        -- B = B - S[2*i+1] 
        "0000000100100111", "0100100000000011",         -- SUB R9, R9, R7
 
        -- B = B >>> A 
        -- initialize R12 with B
        "0000010100101100", "0000000000000000",         -- ADDI R12, R9, 0 
        -- R13 stores A[4:0] - 32 
        "0000110100001101", "0000000000011111",         -- ANDI R13, R8, 31 
        "0000100110101101", "0000000000100000",         -- SUBI R13, R13, 32
        -- R12 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R12 left shift b y 1
        "0000000110001100", "0110000000000001",         -- ADD R12, R12, R12
        -- R13 = R13 + 1 
        "0000010110101101", "0000000000000001",         -- ADDI R13, R13, 1
        -- R12 loop wihle R13 < 0 
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3         
        -- initialize R11 with B
        "0000010100101011", "0000000000000000",         -- ADDI R11, R9, 0
        -- R13 stores A[4:0 ]
        "0000110100001101", "0000000000011111",         -- ANDI R13, R8, 31
        -- R11 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R11 right shift by 1
        "0001010101101011", "0000000000000001",         -- SHR R11, R11, 1 
        -- R13 = R13 -1 
        "0000100110101101", "0000000000000001",         -- SUBI R13, R13, 1 
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3
        -- B = R11 or R12 
        "0000000101101100", "0100100000000111",         -- OR R9, R11, R12 
        -- R11 stores A nor  B
        "0000000100001001", "0101100000001001",         -- NOR R11, R8, R9 
        -- R12 stores A and  B
        "0000000100001001", "0110000000000101",         -- AND R12, R8, R9 

        -- B = A xor B = (A nor B) nor (A and B) 
        "0000000101101100", "0100100000001001",         -- NOR R9, R11, R12 
        -- A = A - S[2*i] 
        "0000000100000110", "0100000000000011",         -- SUB R8, R8, R6 
        -- A = A >>> B 
        -- initialize R12 with A
        "0000010100001100", "0000000000000000",         -- ADDI R12, R8, 0 
        -- R13 stores B[4:0] -32
        "0000110100101101", "0000000000011111",         -- ANDI R13, R9, 31 
        "0000100110101101", "0000000000100000",         -- SUBI R13, R13, 32
        -- R12 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R12 left shift b y 1
        "0000000110001100", "0110000000000001",         -- ADD R12, R12, R12 
        -- R13 = R13 + 1 
        "0000010110101101", "0000000000000001",         -- ADDI R13, R13, 1 
        -- R12 loop wihle R13 < 0
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3 
        -- initialize R11 with A
        "0000010100001011", "0000000000000000",         -- ADDI R11, R8, 0 
        -- R13 stores B[4:0]
        "0000110100101101", "0000000000011111",         -- ANDI R13, R9, 31 
        -- R11 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R11 right shift by 1
        "0001010101101011", "0000000000000001",         -- SHR R11, R11, 1 
        -- R13 = R13 -1 
        "0000100110101101", "0000000000000001",         -- SUBI R13, R13, 1
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3
        "0000000101101100", "0100000000000111",         -- OR R8, R11, R12
        -- R11 stores A nor B
        "0000000100001001", "0101100000001001",         -- NOR R11, R8, R9 
        -- R12 stores A and B
        "0000000100001001", "0110000000000101",         -- AND R12, R8, R9 
        -- A = A xor B = (A nor B) nor (A and B) 
        "0000000101101100", "0100000000001001",         -- NOR R8, R11, R12 
        "0010110000100011", "1111111111010100",         -- BNE R3, R1, -44
        -- R14 = S[0] 
        "0001110000001110", "0000000000000000",         -- LW R14, 0(R0) 
        -- R15 = S[1] 
        "0001110000001111", "0000000000000010",         -- LW R15, 2(R0) 
        -- B = B - S[1] 
        "0000000100101111", "0100100000000011",         -- SUB R9, R9, R15 
        -- A = A - S[0] 
        "0000000100001110", "0100000000000011",         -- SUB R8, R8, R14  
        -- store decrypted A to Mem[52]
        "0010000000001000", "0000000000111000",         -- SW R8, 56(R0) 
        -- store decrypted B to Mem[54]
        "0010000000001001", "0000000000111010",         -- SW R9, 58(R0) 
 
        -- halt 
        "1111110000000000", "0000000000000000",         -- HAL
        others => x"0000"
    );

    -- RC5 key expansion
    constant instr_key : mem := (
        -- initialize part
        "0000000000000001", "0000000000000011",         -- SUB R0, R0, R1 
        "0000010000000100", "0000000000011010",         -- ADDI R4, R0, 26
        "0000010000000101", "0000000000000100",         -- ADDI R5, R0, 4 
        "0000010000000110", "0000000001001110",         -- ADDI R6, R0, 78

        -- L is initialized in data memory based on user input  

        -- initialize S
        -- initialize R1 to be 0
        "0000000000100001", "0000100000000011",         -- SUB R1, R1, R1
        "0001110000000111", "0000000001000100",         -- LW R7, 68(R0)               // R7 <= Mem[68] 0xb7e15163 (magic number P)
        "0010000000000111", "0000000000000000",         -- SW R7, 0(R0)                // Mem[0] <= R7
        "0001110000000111", "0000000001000110",         -- LW R7, 70(R0)               // R7 <= Mem[70] 0xb7e15163 (magic number P)
        "0000010000100001", "0000000000000001",         -- ADDI R1, R1, 1              // R1 <= R1 + 1 (i <= i + 1)
        "0000000000100001", "0100000000000001",         -- ADD R8, R1, R1              // R8 <= R1 << 1 (S loop begin)
        "0001110100001010", "1111111111111110",         -- LW R10, -2(R8)              // R10 <= Mem[R8 - 2] (R10 <= S[i-1])
        "0000000101000111", "0101100000000001",         -- ADD R11, R10, R7            // R11 <= R10 + R7 (R11 <= S[i-1] + Q)
        "0010000100001011", "0000000000000000",         -- SW R11, 0(R8)               // Mem[R8] <= R11 (S[i] <= R11)
        "0000010000100001", "0000000000000001",         -- ADDI R1, R1, 1              // R1 <= R1 + 1 (i <= i + 1)
        "0010110000100100", "1111111111111010",         -- BNE R1, R4, -6              // if R1 != R4, jump to PC + 2 - 12 (S loop end)

        -- mix key into S
        "0000000000100001", "0000100000000011",         -- SUB R1, R1, R1              // R1 <= 0 (i <= 0)
        "0000000001000010", "0001000000000011",         -- SUB R2, R2, R2              // R2 <= 0 (j <= 0)
        "0000000001100011", "0001100000000011",         -- SUB R3, R3, R3              // R3 <= 0 (k <= 0)
        "0000000101001010", "0101000000000011",         -- SUB R10, R10, R10           // R10 <= 0 (A <= 0)
        "0000000101101011", "0101100000000011",         -- SUB R11, R11, R11           // R11 <= 0 (B <= 0)
        -- mix loop begin
        "0000000000100001", "0100000000000001",         -- ADD R8, R1, R1              // R8 <= R1 << 1
        "0000000001000010", "0100100000000001",         -- ADD R9, R2, R2              // R9 <= R2 << 1
        "0000010100101001", "0000000000111100",         -- ADDI R9, R9, 60             // R9 <= R9 + 60
        "0001110100001100", "0000000000000000",         -- LW R12, 0(R8)               // R12 <= Mem[R8] (R12 <= S[i])
        "0001110100101101", "0000000000000000",         -- LW R13, 0(R9)               // R13 <= Mem[R9] (R13 <= L[j])
        -- A <= S[i] + (A + B)
        "0000000101001011", "1000000000000001",         -- ADD R16, R10, R11           // R16 <= R10 + R11
        "0000000110010000", "0101000000000001",         -- ADD R10, R12, R16           // R10 <= R12 + R16
        -- A <= A <<< 3
        "0000010000010000", "0000000000011101",         -- ADDI R16, R0, 29            // R16 <= 29 (loop cycles)
        "0000010101001110", "0000000000000000",         -- ADDI R14, R10, 0            // R14 <= R10 (copy A to R14)
        "0000101000010000", "0000000000000001",         -- SUBI R16, R16, 1            // R16 <= R16 - 1 (R14 loop begin)
        "0001010111001110", "0000000000000001",         -- SHR R14, R14, 1             // R14 <= R14 >> 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R14 loop end)
        "0000010000010000", "0000000000000011",         -- ADDI R16, R0, 3             // R16 <= 3 (loop cycles)
        "0000010101001111", "0000000000000000",         -- ADDI R15, R10, 0            // R15 <= R10 (copy A to R15)
        "0000101000010000", "0000000000000001",         -- SUBI R16, R16, 1            // R16 <= R16 - 1 (R15 loop begin)
        "0000000111101111", "0111100000000001",         -- ADD R15, R15, R15           // R15 <= R15 << 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R15 loop end)
        "0000000111001111", "0101000000000111",         -- OR R10, R14, R15            // R10 <= R14 | R15
        "0010000100001010", "0000000000000000",         -- SW R10, 0(R8)               // Mem[R8] <= R10 (S[i] <= A)
        -- R16 <= (A + B)
        "0000000101001011", "0111100000000001",         -- ADD R15, R10, R11           // R15 <= R10 + R11
        -- B <= L[j] + (A + B)
        "0000000110101111", "0101100000000001",         -- ADD R11, R13, R15           // R11 <= R13 + R15
        -- B <<< (A + B)
        "0000110111110000", "0000000000011111",         -- ANDI R16, R15, 31           // R16 <= R15 & 0x0000001f
        "0000101000010000", "0000000000100000",         -- SUBI R16, R16, 32           // R16 <= R16 - 32
        "0000010101101110", "0000000000000000",         -- ADDI R14, R11, 0            // R14 <= R11 (copy B to R14)
        "0010101000000000", "0000000000000011",         -- BEQ R16, R0, 3              // if R16 = R0, jump to PC + 2 + 6 (R14 loop begin)
        "0000011000010000", "0000000000000001",         -- ADDI R16, R16, 1            // R16 <= R16 + 1
        "0001010111001110", "0000000000000001",         -- SHR R14, R14, 1             // R14 <= R14 >> 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R14 loop end)
        "0000110111110000", "0000000000011111",         -- ANDI R16, R15, 31           // R16 <= R15 & 0x0000001f
        "0000010101101111", "0000000000000000",         -- ADDI R15, R11, 0            // R15 <= R11 (copy B to R15)
        "0010101000000000", "0000000000000011",         -- BEQ R16, R0, 3              // if R16 = R0, jump to PC + 2 + 6 (R15 loop begin)
        "0000101000010000", "0000000000000001",         -- SUBI R16, R16, 1            // R16 <= R16 - 1
        "0000000111101111", "0111100000000001",         -- ADD R15, R15, R15           // R15 <= R15 << 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R15 loop end)
        "0000000111001111", "0101100000000111",         -- OR R11, R14, R15            // R11 <= R14 | R15
        "0010000100101011", "0000000000000000",         -- SW R11, 0(R9)               // Mem[R9] <= R11 (L[j] <= B)
        -- afterthought
        "0000010000100001", "0000000000000001",         -- ADDI R1, R1, 1              // R1 <= R1 + 1 (i <= i + 1)
        "0010110000100100", "0000000000000001",         -- BNE R1, R4, 1               // if R1 != R4, jump to PC + 2 + 2 (if i == 4)
        "0000000000100001", "0000100000000011",         -- SUB R1, R1, R1              // R1 <= 0 (then i <= 0)
        "0000010001000010", "0000000000000001",         -- ADDI R2, R2, 1              // R2 <= R2 + 1 (j <= j + 1)
        "0010110001000101", "0000000000000001",         -- BNE R2, R5, 1               // if R2 != R5, jump to PC + 2 + 2 (if j == 4)
        "0000000001000010", "0001000000000011",         -- SUB R2, R2, R2              // R2 <= 0 (then j <= 0)
        "0000010001100011", "0000000000000001",         -- ADDI R3, R3, 1              // R3 <= R3 + 1 (k <= k + 1)
        "0010110001100110", "1111111111010100",         -- BNE R3, R6, -44             // mix loop end

        -- clear L
        "0000010000000001", "0000000000111100",        -- ADDI R1, R0, 60             // R1 <= 60 (address of L[0])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0
        "0000010000100001", "0000000000000010",        -- ADDI R1, R1, 2              // R1 <= R1 + 2 (find address of L[1])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0
        "0000010000100001", "0000000000000010",        -- ADDI R1, R1, 2              // R1 <= R1 + 2 (find address of L[2])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0
        "0000010000100001", "0000000000000010",        -- ADDI R1, R1, 2              // R1 <= R1 + 2 (find address of L[3])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0

        "1111110000000000", "0000000000000000",         -- HAL 
        others => x"0000"
    );

    -- RC5
    constant instr_rc5 : mem := (
        -- key expansion
        -- initialize part
        "0000000000000001", "0000000000000011",         -- SUB R0, R0, R1 
        "0000010000000100", "0000000000011010",         -- ADDI R4, R0, 26
        "0000010000000101", "0000000000000100",         -- ADDI R5, R0, 4 
        "0000010000000110", "0000000001001110",         -- ADDI R6, R0, 78

        -- L is initialized in data memory based on user input  

        -- initialize S
        -- initialize R1 to be 0
        "0000000000100001", "0000100000000011",         -- SUB R1, R1, R1
        "0001110000000111", "0000000001000100",         -- LW R7, 68(R0)               // R7 <= Mem[68] 0xb7e15163 (magic number P)
        "0010000000000111", "0000000000000000",         -- SW R7, 0(R0)                // Mem[0] <= R7
        "0001110000000111", "0000000001000110",         -- LW R7, 70(R0)               // R7 <= Mem[70] 0xb7e15163 (magic number P)
        "0000010000100001", "0000000000000001",         -- ADDI R1, R1, 1              // R1 <= R1 + 1 (i <= i + 1)
        "0000000000100001", "0100000000000001",         -- ADD R8, R1, R1              // R8 <= R1 << 1 (S loop begin)
        "0001110100001010", "1111111111111110",         -- LW R10, -2(R8)              // R10 <= Mem[R8 - 2] (R10 <= S[i-1])
        "0000000101000111", "0101100000000001",         -- ADD R11, R10, R7            // R11 <= R10 + R7 (R11 <= S[i-1] + Q)
        "0010000100001011", "0000000000000000",         -- SW R11, 0(R8)               // Mem[R8] <= R11 (S[i] <= R11)
        "0000010000100001", "0000000000000001",         -- ADDI R1, R1, 1              // R1 <= R1 + 1 (i <= i + 1)
        "0010110000100100", "1111111111111010",         -- BNE R1, R4, -6              // if R1 != R4, jump to PC + 2 - 12 (S loop end)

        -- mix key into S
        "0000000000100001", "0000100000000011",         -- SUB R1, R1, R1              // R1 <= 0 (i <= 0)
        "0000000001000010", "0001000000000011",         -- SUB R2, R2, R2              // R2 <= 0 (j <= 0)
        "0000000001100011", "0001100000000011",         -- SUB R3, R3, R3              // R3 <= 0 (k <= 0)
        "0000000101001010", "0101000000000011",         -- SUB R10, R10, R10           // R10 <= 0 (A <= 0)
        "0000000101101011", "0101100000000011",         -- SUB R11, R11, R11           // R11 <= 0 (B <= 0)
        -- mix loop begin
        "0000000000100001", "0100000000000001",         -- ADD R8, R1, R1              // R8 <= R1 << 1
        "0000000001000010", "0100100000000001",         -- ADD R9, R2, R2              // R9 <= R2 << 1
        "0000010100101001", "0000000000111100",         -- ADDI R9, R9, 60             // R9 <= R9 + 60
        "0001110100001100", "0000000000000000",         -- LW R12, 0(R8)               // R12 <= Mem[R8] (R12 <= S[i])
        "0001110100101101", "0000000000000000",         -- LW R13, 0(R9)               // R13 <= Mem[R9] (R13 <= L[j])
        -- A <= S[i] + (A + B)
        "0000000101001011", "1000000000000001",         -- ADD R16, R10, R11           // R16 <= R10 + R11
        "0000000110010000", "0101000000000001",         -- ADD R10, R12, R16           // R10 <= R12 + R16
        -- A <= A <<< 3
        "0000010000010000", "0000000000011101",         -- ADDI R16, R0, 29            // R16 <= 29 (loop cycles)
        "0000010101001110", "0000000000000000",         -- ADDI R14, R10, 0            // R14 <= R10 (copy A to R14)
        "0000101000010000", "0000000000000001",         -- SUBI R16, R16, 1            // R16 <= R16 - 1 (R14 loop begin)
        "0001010111001110", "0000000000000001",         -- SHR R14, R14, 1             // R14 <= R14 >> 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R14 loop end)
        "0000010000010000", "0000000000000011",         -- ADDI R16, R0, 3             // R16 <= 3 (loop cycles)
        "0000010101001111", "0000000000000000",         -- ADDI R15, R10, 0            // R15 <= R10 (copy A to R15)
        "0000101000010000", "0000000000000001",         -- SUBI R16, R16, 1            // R16 <= R16 - 1 (R15 loop begin)
        "0000000111101111", "0111100000000001",         -- ADD R15, R15, R15           // R15 <= R15 << 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R15 loop end)
        "0000000111001111", "0101000000000111",         -- OR R10, R14, R15            // R10 <= R14 | R15
        "0010000100001010", "0000000000000000",         -- SW R10, 0(R8)               // Mem[R8] <= R10 (S[i] <= A)
        -- R16 <= (A + B)
        "0000000101001011", "0111100000000001",         -- ADD R15, R10, R11           // R15 <= R10 + R11
        -- B <= L[j] + (A + B)
        "0000000110101111", "0101100000000001",         -- ADD R11, R13, R15           // R11 <= R13 + R15
        -- B <<< (A + B)
        "0000110111110000", "0000000000011111",         -- ANDI R16, R15, 31           // R16 <= R15 & 0x0000001f
        "0000101000010000", "0000000000100000",         -- SUBI R16, R16, 32           // R16 <= R16 - 32
        "0000010101101110", "0000000000000000",         -- ADDI R14, R11, 0            // R14 <= R11 (copy B to R14)
        "0010101000000000", "0000000000000011",         -- BEQ R16, R0, 3              // if R16 = R0, jump to PC + 2 + 6 (R14 loop begin)
        "0000011000010000", "0000000000000001",         -- ADDI R16, R16, 1            // R16 <= R16 + 1
        "0001010111001110", "0000000000000001",         -- SHR R14, R14, 1             // R14 <= R14 >> 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R14 loop end)
        "0000110111110000", "0000000000011111",         -- ANDI R16, R15, 31           // R16 <= R15 & 0x0000001f
        "0000010101101111", "0000000000000000",         -- ADDI R15, R11, 0            // R15 <= R11 (copy B to R15)
        "0010101000000000", "0000000000000011",         -- BEQ R16, R0, 3              // if R16 = R0, jump to PC + 2 + 6 (R15 loop begin)
        "0000101000010000", "0000000000000001",         -- SUBI R16, R16, 1            // R16 <= R16 - 1
        "0000000111101111", "0111100000000001",         -- ADD R15, R15, R15           // R15 <= R15 << 1
        "0010111000000000", "1111111111111101",         -- BNE R16, R0, -3             // if R16 != R0, jump to PC + 2 - 6 (R15 loop end)
        "0000000111001111", "0101100000000111",         -- OR R11, R14, R15            // R11 <= R14 | R15
        "0010000100101011", "0000000000000000",         -- SW R11, 0(R9)               // Mem[R9] <= R11 (L[j] <= B)
        -- afterthought
        "0000010000100001", "0000000000000001",         -- ADDI R1, R1, 1              // R1 <= R1 + 1 (i <= i + 1)
        "0010110000100100", "0000000000000001",         -- BNE R1, R4, 1               // if R1 != R4, jump to PC + 2 + 2 (if i == 4)
        "0000000000100001", "0000100000000011",         -- SUB R1, R1, R1              // R1 <= 0 (then i <= 0)
        "0000010001000010", "0000000000000001",         -- ADDI R2, R2, 1              // R2 <= R2 + 1 (j <= j + 1)
        "0010110001000101", "0000000000000001",         -- BNE R2, R5, 1               // if R2 != R5, jump to PC + 2 + 2 (if j == 4)
        "0000000001000010", "0001000000000011",         -- SUB R2, R2, R2              // R2 <= 0 (then j <= 0)
        "0000010001100011", "0000000000000001",         -- ADDI R3, R3, 1              // R3 <= R3 + 1 (k <= k + 1)
        "0010110001100110", "1111111111010100",         -- BNE R3, R6, -44             // mix loop end

        -- clear L
        "0000010000000001", "0000000000111100",        -- ADDI R1, R0, 60             // R1 <= 60 (address of L[0])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0
        "0000010000100001", "0000000000000010",        -- ADDI R1, R1, 2              // R1 <= R1 + 2 (find address of L[1])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0
        "0000010000100001", "0000000000000010",        -- ADDI R1, R1, 2              // R1 <= R1 + 2 (find address of L[2])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0
        "0000010000100001", "0000000000000010",        -- ADDI R1, R1, 2              // R1 <= R1 + 2 (find address of L[3])
        "0010000000100000", "0000000000000000",        -- SW R0, 0(R1)                // Mem[R1] <= R0

        -- RC5 decryption
        -- initialize part
        -- initialize R0 to 0
        "0000000000000000", "0000000000000011",         -- SUB R0, R0, R0
        -- R3 stores 13 
        "0000010000000011", "0000000000001101",         -- ADDI R3, R0, 13
        -- load A 
        "0001110000001000", "0000000000110100",         -- LW R8, 52(R0)
        -- load B 
        "0001110000001001", "0000000000110110",         -- LW R9, 54(R0)
        -- set R1 as 1 
        "0000010000000001", "0000000000000001",         -- ADDI R1, R0, 1
 
        -- decryption loop begins
        -- R3 = R3 -1 
        "0000100001100011", "0000000000000001",         -- SUBI R3, R3, 1
        -- R4 stores 2*i 
        "0000000001100011", "0010000000000001",         -- ADD R4, R3, R3
        -- R5 stores 2*i+1 
        "0000010010000101", "0000000000000001",         -- ADDI R5, R4, 1 
 
        -- R4 and R5 multiplied by 2 because 16-bit addressable
        "0000000010000100", "0010000000000001",         -- ADD R4, R4, R4
        "0000000010100101", "0010100000000001",         -- ADD R5, R5, R5
        -- R6 stores S[2*i] 
        "0001110010000110", "0000000000000000",         -- LW R6, 0(R4)
        -- R7 stores S[2*i+1]
        "0001110010100111", "0000000000000000",         -- LW R7, 0(R5)
        -- B = B - S[2*i+1] 
        "0000000100100111", "0100100000000011",         -- SUB R9, R9, R7
 
        -- B = B >>> A 
        -- initialize R12 with B
        "0000010100101100", "0000000000000000",         -- ADDI R12, R9, 0 
        -- R13 stores A[4:0] - 32 
        "0000110100001101", "0000000000011111",         -- ANDI R13, R8, 31 
        "0000100110101101", "0000000000100000",         -- SUBI R13, R13, 32
        -- R12 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R12 left shift by 1
        "0000000110001100", "0110000000000001",         -- ADD R12, R12, R12
        -- R13 = R13 + 1 
        "0000010110101101", "0000000000000001",         -- ADDI R13, R13, 1
        -- R12 loop wihle R13 < 0 
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3         
        -- initialize R11 with B
        "0000010100101011", "0000000000000000",         -- ADDI R11, R9, 0
        -- R13 stores A[4:0]
        "0000110100001101", "0000000000011111",         -- ANDI R13, R8, 31
        -- R11 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R11 right shift by 1
        "0001010101101011", "0000000000000001",         -- SHR R11, R11, 1 
        -- R13 = R13 -1 
        "0000100110101101", "0000000000000001",         -- SUBI R13, R13, 1 
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3
        -- B = R11 or R12 
        "0000000101101100", "0100100000000111",         -- OR R9, R11, R12 
        -- R11 stores A nor B
        "0000000100001001", "0101100000001001",         -- NOR R11, R8, R9 
        -- R12 stores A and B
        "0000000100001001", "0110000000000101",         -- AND R12, R8, R9 

        -- B = A xor B = (A nor B) nor (A and B) 
        "0000000101101100", "0100100000001001",         -- NOR R9, R11, R12 
        -- A = A - S[2*i] 
        "0000000100000110", "0100000000000011",         -- SUB R8, R8, R6 
        -- A = A >>> B 
        -- initialize R12 with A
        "0000010100001100", "0000000000000000",         -- ADDI R12, R8, 0 
        -- R13 stores B[4:0] -32
        "0000110100101101", "0000000000011111",         -- ANDI R13, R9, 31 
        "0000100110101101", "0000000000100000",         -- SUBI R13, R13, 32
        -- R12 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R12 left shift by 1
        "0000000110001100", "0110000000000001",         -- ADD R12, R12, R12 
        -- R13 = R13 + 1 
        "0000010110101101", "0000000000000001",         -- ADDI R13, R13, 1 
        -- R12 loop wihle R13 < 0
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3 
        -- initialize R11 with A
        "0000010100001011", "0000000000000000",         -- ADDI R11, R8, 0 
        -- R13 stores B[4:0]
        "0000110100101101", "0000000000011111",         -- ANDI R13, R9, 31 
        -- R11 loop begins 
        "0010100000001101", "0000000000000011",         -- BEQ R13, R0, 3
        -- R11 right shift by 1
        "0001010101101011", "0000000000000001",         -- SHR R11, R11, 1 
        -- R13 = R13 -1 
        "0000100110101101", "0000000000000001",         -- SUBI R13, R13, 1
        "0010110000001101", "1111111111111101",         -- BNE R13, R0, -3
        "0000000101101100", "0100000000000111",         -- OR R8, R11, R12
        -- R11 stores A nor B
        "0000000100001001", "0101100000001001",         -- NOR R11, R8, R9 
        -- R12 stores A and B
        "0000000100001001", "0110000000000101",         -- AND R12, R8, R9 
        -- A = A xor B = (A nor B) nor (A and B) 
        "0000000101101100", "0100000000001001",         -- NOR R8, R11, R12 
        "0010110000100011", "1111111111010100",         -- BNE R3, R1, -44
        -- R14 = S[0] 
        "0001110000001110", "0000000000000000",         -- LW R14, 0(R0) 
        -- R15 = S[1] 
        "0001110000001111", "0000000000000010",         -- LW R15, 2(R0) 
        -- B = B - S[1] 
        "0000000100101111", "0100100000000011",         -- SUB R9, R9, R15 
        -- A = A - S[0] 
        "0000000100001110", "0100000000000011",         -- SUB R8, R8, R14  
        -- store decrypted A to Mem[52]
        "0010000000001000", "0000000000111000",         -- SW R8, 56(R0) 
        -- store decrypted B to Mem[54]
        "0010000000001001", "0000000000111010",         -- SW R9, 58(R0) 
 
        -- halt 
        "1111110000000000", "0000000000000000",         -- HAL
        others => x"0000"
    );
        
end header;