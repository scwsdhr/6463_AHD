library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity instruction_memory is
	port (		
		clr	: in STD_LOGIC;
		A : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		RD : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
end instruction_memory;

architecture Behavioral of instruction_memory is
	
	constant DATA_BITS : INTEGER := 32;			-- number of bits per word
	constant DEPTH     : INTEGER := 256;		-- number of entries
	
	type rom is array (0 to DEPTH - 1) of STD_LOGIC_VECTOR(DATA_BITS - 1 downto 0);
	signal inst_mem : rom := (x"00000000",	
        "00000100000000110000000000000100",
        "00000100000000010000000000000001",
        "00001000011000110000000000000001",
        "00011100011000100000000000000000",
        "00100000011000100000000000001010",
        "00101100000000111111111111111100",
        "00011100000000100000000000001000",
        "00100000000000100000000000001110",
        "00011100000001000000000000001001",
        "00000100000001110000000000011011",
        "00000000100000100001000000010000",
        "00100000001000100000000000001110",
        "00000100001000010000000000000001",
        "00101100111000011111111111111100",
        "00000100000000010000000000000000",
        "00000100001000100000000000000000",
        "00000100001000110000000000000000",
        "00000100001001000000000000000000",
        "00000100001001010000000000000000",
        "00000100000010000000000000000100",
        "00000100000010010000000001001110",
        "00000100000100000000000000011010",
        "00011100001001100000000000001110",
        "00000000100000110001100000010000",
        "00000000110000110001100000010000",
        "00000100000010110000000000000011",
        "00100000000000110000000000110000",
        "00100000000010110000000000110001",
        "00000101011010111111111111111101",
        "00011100000010100000000000101111",
        "00011100000010110000000000110000",
        "00011100000011000000000000110001",
        "00000001010011000110100000010010",
        "00101000000011010000000000001001",
        "00001001101011100000000000100000",
        "00011100000011110000000000110000",
        "00010101011010110000000000000001",
        "00001001101011010000000000000001",
        "00101100000011011111111111111101",
        "00011001111011110000000000000001",
        "00000101110011100000000000000001",
        "00101100000011101111111111111101",
        "00000001111010110101100000010011",
        "00100000001010110000000000001110",
        "00000001011000000001100000010000",
        "00011100010001100000000000001010",
        "00000100100001000000000000000000",
        "00000000100000111010000000010000",
        "00000000110101000010000000010000",
        "00100000000001000000000000110000",
        "00100000000101000000000000110001",
        "00011100000010100000000000101111",
        "00011100000010110000000000110000",
        "00011100000011000000000000110001",
        "00000001010011000110100000010010",
        "00101000000011010000000000001001",
        "00001001101011100000000000100000",
        "00011100000011110000000000110000",
        "00010101011010110000000000000001",
        "00001001101011010000000000000001",
        "00101100000011011111111111111101",
        "00011001111011110000000000000001",
        "00000101110011100000000000000001",
        "00101100000011101111111111111101",
        "00000001111010110101100000010011",
        "00100000010010110000000000001010",
        "00000001011000000010000000010000",
        "00000100001000010000000000000001",
        "00000100010000100000000000000001",
        "00101110000000010000000000000001",
        "00000100000000010000000000000000",
        "00101101000000100000000000000001",
        "00000100000000100000000000000000",
        "00000100101001010000000000000001",
        "00101101001001011111111111001011",
        "00000100000000010000000000000000",
        "00011100001000100000000000001110",
        "00011100001000110000000000101011",
        "00000000011000100001100000010000",
        "00000100001000010000000000000001",
        "00011100001001000000000000001110",
        "00011100001001010000000000101011",
        "00000000101001000010100000010000",
        "00000100000101000000000000001101",
        "00000100001010000000000000000000",
        "00000000101000110011000000010010",
        "00000000101000110011100000010100",
        "00000000111001100011100000010100",
        "00100000000001110000000000110000",
        "00100000000001010000000000110001",
        "00011100000010100000000000101111",
        "00011100000010110000000000110000",
        "00011100000011000000000000110001",
        "00000001010011000110100000010010",
        "00101000000011010000000000001001",
        "00001001101011100000000000100000",
        "00011100000011110000000000110000",
        "00010101011010110000000000000001",
        "00001001101011010000000000000001",
        "00101100000011011111111111111101",
        "00011001111011110000000000000001",
        "00000101110011100000000000000001",
        "00101100000011101111111111111101",
        "00000001111010110101100000010011",
        "00000001000010000100000000010000",
        "00011101000010010000000000001110",
        "00000001001010110001100000010000",
        "00000100011000110000000000000000",
        "00000000101000110011000000010010",
        "00000000101000110011100000010100",
        "00000000111001100011100000010100",
        "00100000000001110000000000110000",
        "00100000000000110000000000110001",
        "00011100000010100000000000101111",
        "00011100000010110000000000110000",
        "00011100000011000000000000110001",
        "00000001010011000110100000010010",
        "00101000000011010000000000001001",
        "00001001101011100000000000100000",
        "00011100000011110000000000110000",
        "00010101011010110000000000000001",
        "00001001101011010000000000000001",
        "00101100000011011111111111111101",
        "00011001111011110000000000000001",
        "00000101110011100000000000000001",
        "00101100000011101111111111111101",
        "00000001111010110101100000010011",
        "00000101000010000000000000000001",
        "00011101000010010000000000001110",
        "00000001001010110010100000010000",
        "00000100101001010000000000000000",
        "00000100001000010000000000000001",
        "00101110100000011111111111010010",
        "00000100000000010000000000000000",
        "00100000001000110000000000101101",
        "00000100011000110000000000000000",
        "00000100001000010000000000000001",
        "00100000001001010000000000101101",
        "00000100101001010000000000000000",
        "00000100000000010000000000000000",
        "00011100001000110000000000101101",
        "00000100001000010000000000000001",
        "00011100001001010000000000101101",
        "00000100000100000000000000000001",
        "00000100000000010000000000001100",
        "00000100001000100000000000000000",
        "00000000001000010000100000010000",
        "00000100001000010000000000000001",
        "00011100001001100000000000001110",
        "00000000110001010010100000010001",
        "00100000000001010000000000110000",
        "00100000000000110000000000110001",
        "00011100000010100000000000101111",
        "00011100000010110000000000110000",
        "00011100000011000000000000110001",
        "00000001010011000110100000010010",
        "00101000000011010000000000001001",
        "00001001101011100000000000100000",
        "00011100000011110000000000110000",
        "00011001011010110000000000000001",
        "00001001101011010000000000000001",
        "00101100000011011111111111111101",
        "00010101111011110000000000000001",
        "00000101110011100000000000000001",
        "00101100000011101111111111111101",
        "00000001111010110101100000010011",
        "00000000011010110100000000010010",
        "00000000011010110011100000010100",
        "00000000111010000010100000010100",
        "00001000001000010000000000000001",
        "00011100001001100000000000001110",
        "00000000110000110001100000010001",
        "00100000000000110000000000110000",
        "00100000000001010000000000110001",
        "00011100000010100000000000101111",
        "00011100000010110000000000110000",
        "00011100000011000000000000110001",
        "00000001010011000110100000010010",
        "00101000000011010000000000001001",
        "00001001101011100000000000100000",
        "00011100000011110000000000110000",
        "00011001011010110000000000000001",
        "00001001101011010000000000000001",
        "00101100000011011111111111111101",
        "00010101111011110000000000000001",
        "00000101110011100000000000000001",
        "00101100000011101111111111111101",
        "00000001111010110101100000010011",
        "00000000101010110100000000010010",
        "00000000101010110011100000010100",
        "00000000111010000001100000010100",
        "00001000001000010000000000000001",
        "00101110000000011111111111010010",
        "00011100001001100000000000001110",
        "00000000110001010010100000010001",
        "00001000001000010000000000000001",
        "00011100001001100000000000001110",
        "00000000110000110001100000010001",
        "00100000000000110000000000101011",
        "00000100011000110000000000000000",
        "00100000000001010000000000101100",
        "00000100101001010000000000000000",
        "11111100000000000000000000000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
        x"00000000",x"00000000",x"00000000",x"00000000",x"00000000");

begin

	process(clr)
	begin
		if (clr = '1') then
            null;
 		end if;
	end process;
	
	RD <= inst_mem(conv_integer(A));	
	
end Behavioral;